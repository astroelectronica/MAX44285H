.title KiCad schematic
.include "C:/AE/MAX44285H/_models/C2012C0G2A102J060AA_p.mod"
.include "C:/AE/MAX44285H/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/MAX44285H/_models/max44285.lib"
R3 VCC /LOAD1 {RSNS1}
R4 VCC /LOAD2 {RSNS2}
I2 /LOAD1 0 {LOAD1}
I1 /LOAD2 0 {LOAD2}
R1 /VOCM1 /OUT1 {RLPF1}
XU1 /OUT1 0 C2012C0G2A102J060AA_p
XU2 /OUT2 0 C2012C0G2A102J060AA_p
XU4 VDD 0 C2012X7R2A104K125AA_p
XU3 VCC /LOAD1 /VOCM1 VCC /LOAD2 /VOCM2 VDD 0 MAX44285H
V1 VDD 0 {VSUPPLY}
V2 VCC 0 {VSOURCE}
R2 /VOCM2 /OUT2 {RLPF2}
.end
